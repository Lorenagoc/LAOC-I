library verilog;
use verilog.vl_types.all;
entity FUNC2 is
    port(
        \out\           : out    vl_logic_vector(7 downto 0);
        ctl             : in     vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
end FUNC2;
