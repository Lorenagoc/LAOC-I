library verilog;
use verilog.vl_types.all;
entity B_15 is
    port(
        HAB             : in     vl_logic;
        D               : in     vl_logic;
        Q               : out    vl_logic
    );
end B_15;
